* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT INV_2X OUT IN VDD GND
** N=4 EP=4 IP=0 FDC=2
M0 GND IN OUT GND N_18 L=1.8e-07 W=5.1e-07 AD=4.488e-13 AS=4.386e-13 PD=2.27e-06 PS=2.23e-06 $X=18540 $Y=4710 $D=0
M1 VDD IN OUT VDD P_18 L=1.8e-07 W=5.3e-07 AD=4.24e-13 AS=4.505e-13 PD=2.13e-06 PS=2.23e-06 $X=18540 $Y=10780 $D=1
.ENDS
***************************************
.SUBCKT MUX21 out in1 in2 ctrl GND VDD
** N=7 EP=6 IP=0 FDC=6
M0 out ctrl in2 GND N_18 L=1.8e-07 W=5e-07 AD=3.225e-13 AS=5.675e-13 PD=1.29e-06 PS=2.77e-06 $X=27735 $Y=12070 $D=0
M1 in1 7 out GND N_18 L=1.8e-07 W=5e-07 AD=4.225e-13 AS=3.225e-13 PD=2.19e-06 PS=1.29e-06 $X=29205 $Y=12070 $D=0
M2 GND ctrl 7 GND N_18 L=1.8e-07 W=5e-07 AD=4.55e-13 AS=4.7e-13 PD=2.32e-06 PS=2.38e-06 $X=31550 $Y=12070 $D=0
M3 out ctrl in1 VDD P_18 L=1.8e-07 W=5.7e-07 AD=3.6765e-13 AS=6.2985e-13 PD=1.29e-06 PS=2.78e-06 $X=27735 $Y=18100 $D=1
M4 in2 7 out VDD P_18 L=1.8e-07 W=5.7e-07 AD=4.7025e-13 AS=3.6765e-13 PD=2.22e-06 PS=1.29e-06 $X=29205 $Y=18100 $D=1
M5 VDD ctrl 7 VDD P_18 L=1.8e-07 W=5.7e-07 AD=5.244e-13 AS=5.358e-13 PD=2.41e-06 PS=2.45e-06 $X=31550 $Y=18100 $D=1
.ENDS
***************************************
.SUBCKT FA VDD b a GND c_in c_out sum
** N=12 EP=7 IP=38 FDC=34
X0 8 a VDD GND INV_2X $T=4350 -16930 0 0 $X=21530 $Y=-13700
X1 11 12 VDD GND INV_2X $T=17620 -16930 0 0 $X=34800 $Y=-13700
X2 9 GND a b GND VDD MUX21 $T=-4470 -36240 0 0 $X=21620 $Y=-26110
X3 12 a 8 b GND VDD MUX21 $T=-50 -24340 0 0 $X=26040 $Y=-14210
X4 10 a VDD b GND VDD MUX21 $T=4430 -36240 0 0 $X=30520 $Y=-26110
X5 c_out 9 10 c_in GND VDD MUX21 $T=13150 -36240 0 0 $X=39240 $Y=-26110
X6 sum 12 11 c_in GND VDD MUX21 $T=13170 -24340 0 0 $X=39260 $Y=-14210
.ENDS
***************************************
.SUBCKT ADDER3 VDD A0 GND B1 A1 CIN A2 S2 COUT S1 SO B0 B2
** N=25 EP=13 IP=66 FDC=228
X0 S2 17 13 CIN GND VDD MUX21 $T=107500 -40190 0 180 $X=74310 $Y=-60790
X1 COUT 14 12 CIN GND VDD MUX21 $T=107500 -28220 0 180 $X=74310 $Y=-48820
X2 S1 9 4 CIN GND VDD MUX21 $T=48350 -43590 0 0 $X=74440 $Y=-33460
X3 SO 11 8 CIN GND VDD MUX21 $T=48350 -31440 0 0 $X=74440 $Y=-21310
X4 VDD B0 A0 GND VDD 2 8 FA $T=59880 -64460 0 180 $X=11730 $Y=-60720
X5 VDD B0 A0 GND GND 22 11 FA $T=-8520 -7060 0 0 $X=12590 $Y=-33780
X6 VDD B1 A1 GND 2 23 4 FA $T=90680 -64460 0 180 $X=42530 $Y=-60720
X7 VDD B1 A1 GND 22 16 9 FA $T=21800 -7060 0 0 $X=42910 $Y=-33780
X8 VDD B2 A2 GND 23 12 13 FA $T=133150 -64460 0 180 $X=85000 $Y=-60720
X9 VDD B2 A2 GND 16 14 17 FA $T=64750 -7060 0 0 $X=85860 $Y=-33780
.ENDS
***************************************
