* SPICE NETLIST
***************************************

.SUBCKT L POS NEG
.ENDS
***************************************
.SUBCKT INV_2X OUT IN VDD GND
** N=4 EP=4 IP=0 FDC=2
M0 GND IN OUT GND N_18 L=1.8e-07 W=5.1e-07 AD=4.488e-13 AS=4.386e-13 PD=2.27e-06 PS=2.23e-06 $X=18540 $Y=4710 $D=0
M1 VDD IN OUT VDD P_18 L=1.8e-07 W=5.3e-07 AD=4.24e-13 AS=4.505e-13 PD=2.13e-06 PS=2.23e-06 $X=18540 $Y=10780 $D=1
.ENDS
***************************************
.SUBCKT MUX21 out in1 in2 ctrl GND VDD
** N=7 EP=6 IP=0 FDC=6
M0 out ctrl in2 GND N_18 L=1.8e-07 W=5e-07 AD=3.225e-13 AS=5.675e-13 PD=1.29e-06 PS=2.77e-06 $X=27735 $Y=12070 $D=0
M1 in1 7 out GND N_18 L=1.8e-07 W=5e-07 AD=4.225e-13 AS=3.225e-13 PD=2.19e-06 PS=1.29e-06 $X=29205 $Y=12070 $D=0
M2 GND ctrl 7 GND N_18 L=1.8e-07 W=5e-07 AD=4.55e-13 AS=4.7e-13 PD=2.32e-06 PS=2.38e-06 $X=31550 $Y=12070 $D=0
M3 out ctrl in1 VDD P_18 L=1.8e-07 W=5.7e-07 AD=3.6765e-13 AS=6.2985e-13 PD=1.29e-06 PS=2.78e-06 $X=27735 $Y=18100 $D=1
M4 in2 7 out VDD P_18 L=1.8e-07 W=5.7e-07 AD=4.7025e-13 AS=3.6765e-13 PD=2.22e-06 PS=1.29e-06 $X=29205 $Y=18100 $D=1
M5 VDD ctrl 7 VDD P_18 L=1.8e-07 W=5.7e-07 AD=5.244e-13 AS=5.358e-13 PD=2.41e-06 PS=2.45e-06 $X=31550 $Y=18100 $D=1
.ENDS
***************************************
.SUBCKT FA VDD b a GND c_in c_out sum
** N=12 EP=7 IP=38 FDC=34
X0 2 a VDD GND INV_2X $T=4350 -16930 0 0 $X=21530 $Y=-13700
X1 7 8 VDD GND INV_2X $T=17620 -16930 0 0 $X=34800 $Y=-13700
X2 3 GND a b GND VDD MUX21 $T=-4470 -36240 0 0 $X=21620 $Y=-26110
X3 8 a 2 b GND VDD MUX21 $T=-50 -24340 0 0 $X=26040 $Y=-14210
X4 6 a VDD b GND VDD MUX21 $T=4430 -36240 0 0 $X=30520 $Y=-26110
X5 c_out 3 6 c_in GND VDD MUX21 $T=13150 -36240 0 0 $X=39240 $Y=-26110
X6 sum 8 7 c_in GND VDD MUX21 $T=13170 -24340 0 0 $X=39260 $Y=-14210
.ENDS
***************************************
